library verilog;
use verilog.vl_types.all;
entity adder_4bit is
    port(
        a               : in     vl_logic_vector(3 downto 0);
        b               : in     vl_logic_vector(3 downto 0);
        carry_in        : in     vl_logic;
        sum             : out    vl_logic_vector(3 downto 0);
        overflow        : out    vl_logic
    );
end adder_4bit;
