library verilog;
use verilog.vl_types.all;
entity tb_sda_sel is
end tb_sda_sel;
