// $Id: $
// File name:   adder_nbit.sv
// Created:     1/22/2015
// Author:      Parneet Kaur Ahuja
// Lab Section: 01
// Version:     1.0  Initial Design Entry
// Description: n bit adder
`timescale 1ns / 100ps
module adder_nbit
#(
  parameter num = 16
)
(
	input wire [(num - 1):0] a,
	input wire [(num - 1):0] b,
	input wire carry_in,
	output wire [(num - 1):0] sum,
	output wire overflow
);
wire [num:0] carrys;
genvar i;
assign carrys[0] = carry_in;

generate
  for(i = 0; i <= (num - 1); i = i + 1)
  begin
    adder_1bit Ii (.a(a[i]), .b(b[i]), .carry_in(carrys[i]), .sum(sum[i]), .carry_out(carrys[i+1]));
    always @ (a)
  begin
    assert((a[i] == 1'b1) || (a[i] == 1'b0))
  else $error("Input 'a' of component is not a digital logic value");
  end
  always @ (b)
  begin
    assert((b[i] == 1'b1) || (b[i] == 1'b0))
  else $error("Input 'b' of component is not a digital logic value");
  end
  always @ (carry_in)
  begin
    assert((carry_in == 1'b1) || (carry_in == 1'b0))
  else $error("Input 'carry_in' of component is not a digital logic value");
  end
   
    always @(a[i],b[i],carrys[i])
    begin
    #(2) assert(((a[i] +b[i] + carrys[i]) % 2) == sum[i])
    else $error("Output 's' of first 1 bit adder is not correct");
    end
  end
  
endgenerate
assign overflow = carrys[num];
endmodule