library verilog;
use verilog.vl_types.all;
entity flex_counter_NUM_CNT_BITS10_DW01_inc_0 is
    port(
        A               : in     vl_logic_vector(9 downto 0);
        SUM             : out    vl_logic_vector(9 downto 0)
    );
end flex_counter_NUM_CNT_BITS10_DW01_inc_0;
