library verilog;
use verilog.vl_types.all;
entity scl_edge is
    port(
        clk             : in     vl_logic;
        n_rst           : in     vl_logic;
        scl             : in     vl_logic;
        falling_edge_found: out    vl_logic;
        rising_edge_found: out    vl_logic
    );
end scl_edge;
