library verilog;
use verilog.vl_types.all;
entity tb_tx_fifo is
end tb_tx_fifo;
