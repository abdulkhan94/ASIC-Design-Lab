`timescale 1ns / 10ps

module tb_test();

localparam	CLK_PERIOD		= 2.5;

reg clk;
reg n_rst;


always
begin
	clk = 1'b0;
	#(CLK_PERIOD/2.0);
	clk = 1'b1;
	#(CLK_PERIOD/2.0);
end



reg start_byte;
reg stop_byte;

reg master_readdatavalid;
reg master_waitrequest;

test DUT(
	.clk(clk),
	.reset_n(n_rst),
	.stop_byte(stop_byte),
	.start_byte(start_byte),
	.master_readdatavalid(master_readdatavalid),
	.master_waitrequest(master_waitrequest)
);

initial
	begin
	n_rst = 1;
	#(CLK_PERIOD);
	n_rst = 0;
	#(CLK_PERIOD);
	n_rst = 1;
	
	#(CLK_PERIOD);
	start_byte = 1;
	#(4*CLK_PERIOD);
	master_readdatavalid = 1;
	master_waitrequest = 0;
	#(CLK_PERIOD*20);
	

end

endmodule

