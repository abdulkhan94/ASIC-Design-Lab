library verilog;
use verilog.vl_types.all;
entity tb_adder_8bit is
end tb_adder_8bit;
