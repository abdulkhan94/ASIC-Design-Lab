// $Id: $
// File name:   adder_1bit.sv
// Created:     1/27/2015
// Author:      Parneet Kaur Ahuja
// Lab Section: 01
// Version:     1.0  Initial Design Entry
// Description: 1 bit full adder

`timescale 1ns / 100ps
module adder_1bit
(
	input wire  a,
	input wire  b,
	input wire carry_in,
	output wire sum,
	output wire carry_out
);
wire mid1;
wire mid2;
wire mid3;
wire mid4;
wire mid5;

	xor a1 (mid1, a, b);
  xor a2 (sum, mid1, carry_in);
  or a3 (mid2, b, a);
  and a4 (mid3, carry_in, mid2);
  and a5 (mid4, b, a);
  and a6 (mid5, mid4, !carry_in);
  or a7 (carry_out, mid5, mid3);	
  
  always @ (a)
  begin
    assert((a == 1'b1) || (a == 1'b0))
  else $error("Input 'a' of component is not a digital logic value");
  end
  always @ (b)
  begin
    assert((b == 1'b1) || (b == 1'b0))
  else $error("Input 'b' of component is not a digital logic value");
  end
  always @ (carry_in)
  begin
    assert((carry_in == 1'b1) || (carry_in == 1'b0))
  else $error("Input 'carry_in' of component is not a digital logic value");
  end
    
endmodule